module not_gate(
    input wire a,
    output wire out
);
    assign out = ~a;
endmodule
