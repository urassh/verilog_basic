module tb_full_adder;

endmodule
