module not(
    input wire a,
    output wire out;
);
    assign out = ~a;
endmodule
